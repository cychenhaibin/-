library verilog;
use verilog.vl_types.all;
entity m6 is
    port(
        co_34           : out    vl_logic_vector(2 downto 0);
        clk8_34         : in     vl_logic
    );
end m6;
