library verilog;
use verilog.vl_types.all;
entity spead_select_vlg_vec_tst is
end spead_select_vlg_vec_tst;
