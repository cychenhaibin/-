library verilog;
use verilog.vl_types.all;
entity m10_vlg_check_tst is
    port(
        co_34           : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end m10_vlg_check_tst;
