library verilog;
use verilog.vl_types.all;
entity dig_select_34 is
    port(
        q_34            : out    vl_logic_vector(7 downto 0);
        p_34            : in     vl_logic_vector(2 downto 0)
    );
end dig_select_34;
