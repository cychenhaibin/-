library verilog;
use verilog.vl_types.all;
entity counter100_vlg_vec_tst is
end counter100_vlg_vec_tst;
