library verilog;
use verilog.vl_types.all;
entity m10 is
    port(
        q_000           : out    vl_logic_vector(3 downto 0);
        input           : in     vl_logic
    );
end m10;
