library verilog;
use verilog.vl_types.all;
entity dig_select_34_vlg_check_tst is
    port(
        q_34            : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end dig_select_34_vlg_check_tst;
