library verilog;
use verilog.vl_types.all;
entity cnt24_8_vlg_vec_tst is
end cnt24_8_vlg_vec_tst;
