library verilog;
use verilog.vl_types.all;
entity cnt6 is
    port(
        q_000           : out    vl_logic_vector(2 downto 0);
        i_16            : in     vl_logic
    );
end cnt6;
