library verilog;
use verilog.vl_types.all;
entity cnt16_vlg_vec_tst is
end cnt16_vlg_vec_tst;
