library verilog;
use verilog.vl_types.all;
entity demo2_34_vlg_vec_tst is
end demo2_34_vlg_vec_tst;
