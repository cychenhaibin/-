library verilog;
use verilog.vl_types.all;
entity common_clock_vlg_vec_tst is
end common_clock_vlg_vec_tst;
