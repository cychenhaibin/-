library verilog;
use verilog.vl_types.all;
entity m10_vlg_vec_tst is
end m10_vlg_vec_tst;
