library verilog;
use verilog.vl_types.all;
entity tell_time_vlg_vec_tst is
end tell_time_vlg_vec_tst;
