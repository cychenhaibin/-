library verilog;
use verilog.vl_types.all;
entity cnt7_vlg_vec_tst is
end cnt7_vlg_vec_tst;
