library verilog;
use verilog.vl_types.all;
entity m10_vlg_sample_tst is
    port(
        clk_34          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end m10_vlg_sample_tst;
