library verilog;
use verilog.vl_types.all;
entity spead_select_vlg_check_tst is
    port(
        outhz_34        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end spead_select_vlg_check_tst;
