library verilog;
use verilog.vl_types.all;
entity counter60_vlg_vec_tst is
end counter60_vlg_vec_tst;
