library verilog;
use verilog.vl_types.all;
entity cnt60 is
    port(
        q_13            : out    vl_logic;
        clk_60          : in     vl_logic;
        q_12            : out    vl_logic;
        q_100           : out    vl_logic;
        q_101           : out    vl_logic;
        q_10            : out    vl_logic;
        q_11            : out    vl_logic;
        q_103           : out    vl_logic;
        q_102           : out    vl_logic
    );
end cnt60;
