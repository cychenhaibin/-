library verilog;
use verilog.vl_types.all;
entity cnt24_8_vlg_sample_tst is
    port(
        clk_24_8        : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end cnt24_8_vlg_sample_tst;
