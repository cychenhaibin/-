library verilog;
use verilog.vl_types.all;
entity key_debounce_vlg_check_tst is
    port(
        key_out_000     : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end key_debounce_vlg_check_tst;
