library verilog;
use verilog.vl_types.all;
entity bell_music_vlg_check_tst is
    port(
        bell_go         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end bell_music_vlg_check_tst;
