library verilog;
use verilog.vl_types.all;
entity counter24_vlg_vec_tst is
end counter24_vlg_vec_tst;
