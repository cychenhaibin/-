library verilog;
use verilog.vl_types.all;
entity m10_vlg_check_tst is
    port(
        co              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end m10_vlg_check_tst;
