library verilog;
use verilog.vl_types.all;
entity docker_34_vlg_vec_tst is
end docker_34_vlg_vec_tst;
