library verilog;
use verilog.vl_types.all;
entity cnt10_vlg_check_tst is
    port(
        co              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end cnt10_vlg_check_tst;
