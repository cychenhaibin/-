library verilog;
use verilog.vl_types.all;
entity docker_34 is
    port(
        seg_34          : out    vl_logic_vector(6 downto 0);
        d_34            : in     vl_logic_vector(3 downto 0)
    );
end docker_34;
