library verilog;
use verilog.vl_types.all;
entity m10 is
    port(
        co_34           : out    vl_logic_vector(3 downto 0);
        clk_34          : in     vl_logic
    );
end m10;
