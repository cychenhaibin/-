library verilog;
use verilog.vl_types.all;
entity code_select_8_vlg_vec_tst is
end code_select_8_vlg_vec_tst;
