library verilog;
use verilog.vl_types.all;
entity key_debounce_vlg_vec_tst is
end key_debounce_vlg_vec_tst;
