library verilog;
use verilog.vl_types.all;
entity cnt60_vlg_check_tst is
    port(
        q_10            : in     vl_logic;
        q_11            : in     vl_logic;
        q_12            : in     vl_logic;
        q_13            : in     vl_logic;
        q_100           : in     vl_logic;
        q_101           : in     vl_logic;
        q_102           : in     vl_logic;
        q_103           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end cnt60_vlg_check_tst;
