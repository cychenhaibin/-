library verilog;
use verilog.vl_types.all;
entity m6_vlg_vec_tst is
end m6_vlg_vec_tst;
