library verilog;
use verilog.vl_types.all;
entity bell_music_vlg_vec_tst is
end bell_music_vlg_vec_tst;
