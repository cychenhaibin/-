library verilog;
use verilog.vl_types.all;
entity knocker_vlg_vec_tst is
end knocker_vlg_vec_tst;
