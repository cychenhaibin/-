library verilog;
use verilog.vl_types.all;
entity cnt24_34_vlg_sample_tst is
    port(
        clear24_34      : in     vl_logic;
        clk_cnt24_34    : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end cnt24_34_vlg_sample_tst;
