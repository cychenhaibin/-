library verilog;
use verilog.vl_types.all;
entity cnt60_34_vlg_sample_tst is
    port(
        clear60_34      : in     vl_logic;
        clk_cnt60_34    : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end cnt60_34_vlg_sample_tst;
