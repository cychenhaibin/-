library verilog;
use verilog.vl_types.all;
entity knocker_vlg_check_tst is
    port(
        bee_000         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end knocker_vlg_check_tst;
